module lab5_1
    
